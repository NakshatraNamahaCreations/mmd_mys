�PNG

   IHDR         rߔ   sRGB ���  (IDATHŖ�� �YC:Fgp���
]�c���܁k�G�z��"r���ȗ��XB㢩+�~�Њ� �z��~��D-/�IzrI��&uI{��f���sA�&4_� # z>�_�ùk/��3�5'�F�o��A�y@�t��3[SR�ɘ��A��ͻ�'ѻ)��*&I[+q�O8�����Y"{��`1����[�s���: ϸ{1�%@<71�r�å���-8"O�+�EዏtS4�X<y[+��� �G��y��l���5m���J ъQ���[�L�P|m��(��P��,��T��py�    IEND�B`�